package write_fsm_pkg is
	type write_fsm_state_type is ( idl_rdt, cmp_sto, wait_sto);
end package write_fsm_pkg;

--package body write_fsm_pkg is
--
--end package body write_fsm_pkg;

