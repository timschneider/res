package read_fsm_pkg is
	type read_fsm_state_type is ( idl_rdt, cmp_dlv, req0, req1,rd0,rd1, rd1_keep,rd2,rd3,rd4,rd5,rd6,rd7, sync);
end package read_fsm_pkg;

